`ifndef __RISC_INST_CONSTANTS__
    `define __RISC_INST_CONSTANTS__



`define  MEMORY_CODE_START_ADDR      0
`define  MEMORY_CODE_END_ADDR       10
`define  REGFILE_SIZE				32


`endif