
//`include "risc_scoreboard.sv"

`include "risc_test_top.sv"






